module instrMem (
    input wire clk,
    input wire rst,
    input wire [31:0] addr,
    output reg [31:0] data
);
    //reg [31:0] mem [0:(2**32)-1];
    reg [31:0] mem [0:31];

    initial begin
        mem[0]  = 32'b10001100000000010000000000000001;
        mem[1]  = 32'b10001100000000100000000000000010;
        mem[2]  = 32'b10001100000000110000000000000011;
        mem[3]  = 32'b10000000000000000000000000000000;
        mem[4]  = 32'b10000000000000000000000000000000;
        mem[5]  = 32'b00000000001000100000100000100000;
        mem[6]  = 32'b10000000000000000000000000000000;
        mem[7]  = 32'b10000000000000000000000000000000;
        mem[8]  = 32'b10000000000000000000000000000000;
        mem[9]  = 32'b00000000001000110000100000100000;
        mem[10] = 32'b10000000000000000000000000000000;
        mem[11] = 32'b10000000000000000000000000000000;
        mem[12] = 32'b10000000000000000000000000000000;
        mem[13] = 32'b00000000001000010000100000100000;
        mem[14] = 32'b10000000000000000000000000000000;
        mem[15] = 32'b10000000000000000000000000000000;
        mem[16] = 32'b10000000000000000000000000000000;
        mem[17] = 32'b10000000000000000000000000000000;
        mem[18] = 32'b00000000001000000000100000100000;
        mem[19] = 32'b10000000000000000000000000000000;
        mem[20] = 32'b10000000000000000000000000000000;
        mem[21] = 32'b10000000000000000000000000000000;
        mem[22] = 32'b10000000000000000000000000000000;
        mem[23] = 32'b10000000000000000000000000000000;
    end

    always @(*) begin
        data = mem[addr[31:2]];
    end
endmodule
